

 
 
 




window new WaveWindow  -name  "Waves for BMG Example Design"
waveform  using  "Waves for BMG Example Design"

      waveform add -signals /Block_Memory_64x24_tb/status
      waveform add -signals /Block_Memory_64x24_tb/Block_Memory_64x24_synth_inst/bmg_port/CLKA
      waveform add -signals /Block_Memory_64x24_tb/Block_Memory_64x24_synth_inst/bmg_port/ADDRA
      waveform add -signals /Block_Memory_64x24_tb/Block_Memory_64x24_synth_inst/bmg_port/DINA
      waveform add -signals /Block_Memory_64x24_tb/Block_Memory_64x24_synth_inst/bmg_port/WEA
      waveform add -signals /Block_Memory_64x24_tb/Block_Memory_64x24_synth_inst/bmg_port/RSTB
      waveform add -signals /Block_Memory_64x24_tb/Block_Memory_64x24_synth_inst/bmg_port/CLKB
      waveform add -signals /Block_Memory_64x24_tb/Block_Memory_64x24_synth_inst/bmg_port/ADDRB
      waveform add -signals /Block_Memory_64x24_tb/Block_Memory_64x24_synth_inst/bmg_port/DOUTB

console submit -using simulator -wait no "run"
